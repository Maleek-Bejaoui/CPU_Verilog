----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 16.01.2025 10:26:21
-- Design Name: 
-- Module Name: Accu_register - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Accu_register is
    Port (  clk         : in STD_LOGIC;
            ce          : in STD_LOGIC;
            rst         : in STD_LOGIC;
            load_ACCU   : in STD_LOGIC;
            data_in     : in STD_LOGIC_VECTOR (15 downto 0);
            data_out    : out STD_LOGIC_VECTOR (15 downto 0));
end Accu_register;

architecture Behavioral of Accu_register is

begin

    process(rst, clk)
        begin
        if(rst = '1') then
            data_out <= (others => '0');
        elsif(rising_edge(clk)) then
            if(ce = '1') then
                if (load_ACCU = '1') then 
                    data_out <= data_in;
                end if;
            end if;
        end if;
    end process;
    
end Behavioral;
